library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity HYGRO_handler is
--    Port(
    
--    );
end HYGRO_handler;

architecture Behavioral of HYGRO_handler is

begin


end Behavioral;
